module K_value_g_Holder (
 
  output reg [15:0] value
);

 
    initial begin
      value <= 16'hFF00;
    end
  

endmodule


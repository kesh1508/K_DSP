module K_value_b_Holder (
  
  output reg [15:0] value
);

  
   initial begin 
      value <= 16'h00FF;
    
  end

endmodule

